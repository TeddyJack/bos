module ram_control
(
  fsdf
);


endmodule