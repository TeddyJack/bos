module cmd_encoder(
output [7:0] tx_data,
output       tx_valid,
input        tx_ready
);


endmodule